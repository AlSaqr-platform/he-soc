/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */
// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 319;
    const logic [RomSize-1:0][63:0] mem = {
         64'h000000000000000A,
         64'h4645444342413938,
         64'h3736353433323130,
         64'h00000000FF5FF06F,
         64'hDF1FF0EFDBDFF0EF,
         64'hD8DFF0EF00113423,
         64'hFF010113FFDFF06F,
         64'h1050007300E7F663,
         64'h00100793F1402773,
         64'h68858593FFFFF597,
         64'hF1402573E5DFF06F,
         64'h0201011301813083,
         64'h00914503E6DFF0EF,
         64'h00814503F09FF0EF,
         64'h00113C2300810593,
         64'hFE01011300008067,
         64'h0301011301013903,
         64'h0181348302013403,
         64'h02813083FD241EE3,
         64'hEA1FF0EF00914503,
         64'hEA9FF0EFFF84041B,
         64'h00814503F49FF0EF,
         64'h0FF5751300810593,
         64'h0084D533FF800913,
         64'h0380041300050493,
         64'h0211342301213823,
         64'h00913C2302813023,
         64'hFD01011300008067,
         64'h0301011301013903,
         64'h0181348302013403,
         64'h02813083FD241EE3,
         64'hF01FF0EF00914503,
         64'hF09FF0EFFF84041B,
         64'h00814503FA9FF0EF,
         64'h0FF5751300810593,
         64'h0084D53BFF800913,
         64'h0180041300050493,
         64'h0211342301213823,
         64'h00913C2302813023,
         64'hFD01011300008067,
         64'h00F580230007C783,
         64'h00E580A300A787B3,
         64'h0045551300074703,
         64'h00E7873300F57713,
         64'h1507879300000797,
         64'hFE1FF06F00140413,
         64'hF79FF0EF00008067,
         64'h0101011300013403,
         64'h0081308300051A63,
         64'h0004450300050413,
         64'h0011342300813023,
         64'hFF01011300008067,
         64'h00E7882302000713,
         64'h00E78423FC700713,
         64'h00E7862300300713,
         64'h00A782230FF57513,
         64'h00E780230085551B,
         64'h0FF5771300E78623,
         64'hF800071300078223,
         64'h400007B702B5553B,
         64'h0045959B00008067,
         64'h00A70023FE078CE3,
         64'h0207F79301474783,
         64'h4000073700008067,
         64'h020575130147C503,
         64'h400007B700008067,
         64'h0005450300008067,
         64'h00B5002300008067,
         64'h0002806700056283,
         64'h104045370207A223,
         64'h104047B700008067,
         64'h0807A0230C0027B7,
         64'h00F722230C201737,
         64'h000080671807A023,
         64'h0C0027B700F72223,
         64'h0C20373700070C63,
         64'h2607A78300000797,
         64'hF1402773FDDFF06F,
         64'h0C2037B700008067,
         64'hFEE698E328072703,
         64'h0007A68300000717,
         64'h105000730080006F,
         64'h004787930C2017B7,
         64'h02079463F14027F3,
         64'h0000806700000000,
         64'h68746469772D6F69,
         64'h2D67657200746669,
         64'h68732D6765720073,
         64'h747075727265746E,
         64'h6900746E65726170,
         64'h2D74707572726574,
         64'h6E69006465657073,
         64'h2D746E6572727563,
         64'h007665646E2C7663,
         64'h7369720079746972,
         64'h6F6972702D78616D,
         64'h2C76637369720073,
         64'h656D616E2D676572,
         64'h006465646E657478,
         64'h652D737470757272,
         64'h65746E6900736567,
         64'h6E617200656C646E,
         64'h6168700072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h00736C6C65632D74,
         64'h7075727265746E69,
         64'h230074696C70732D,
         64'h626C740065707974,
         64'h2D756D6D00617369,
         64'h2C76637369720079,
         64'h636E657571657266,
         64'h2D6B636F6C630073,
         64'h7574617473007963,
         64'h6E6575716572662D,
         64'h65736162656D6974,
         64'h0067657200657079,
         64'h745F656369766564,
         64'h00687461702D7475,
         64'h6F647473006C6564,
         64'h6F6D00656C626974,
         64'h61706D6F6300736C,
         64'h6C65632D657A6973,
         64'h2300736C6C65632D,
         64'h7373657264646123,
         64'h0900000002000000,
         64'h0200000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000002000000,
         64'h0E01000004000000,
         64'h0300000000100000,
         64'h0000000000000018,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0700000006000000,
         64'h0500000004000000,
         64'h1F01000010000000,
         64'h0300000000007265,
         64'h6D69745F6270612C,
         64'h706C75701B000000,
         64'h0F00000003000000,
         64'h0000303030303030,
         64'h38314072656D6974,
         64'h0100000002000000,
         64'h0400000034010000,
         64'h0400000003000000,
         64'h020000002A010000,
         64'h0400000003000000,
         64'h020000001F010000,
         64'h0400000003000000,
         64'h020000000E010000,
         64'h0400000003000000,
         64'h00C2010000010000,
         64'h0400000003000000,
         64'h80F0FA0262000000,
         64'h0400000003000000,
         64'h0010000000000000,
         64'h0000004000000000,
         64'h4400000010000000,
         64'h0300000000303535,
         64'h3631736E1B000000,
         64'h0800000003000000,
         64'h0000003030303030,
         64'h3030344074726175,
         64'h0100000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000000100000,
         64'h0000000000000000,
         64'h0000000044000000,
         64'h1000000003000000,
         64'hFFFF000001000000,
         64'hC400000008000000,
         64'h0300000000333130,
         64'h2D67756265642C76,
         64'h637369721B000000,
         64'h1000000003000000,
         64'h0000304072656C6C,
         64'h6F72746E6F632D67,
         64'h7562656401000000,
         64'h0200000002000000,
         64'hB500000004000000,
         64'h03000000FF000000,
         64'hF500000004000000,
         64'h0300000007000000,
         64'hE200000004000000,
         64'h0300000000000004,
         64'h000000000000000C,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0900000001000000,
         64'h0B00000001000000,
         64'hC400000010000000,
         64'h03000000A0000000,
         64'h0000000003000000,
         64'h003063696C702C76,
         64'h637369721B000000,
         64'h0C00000003000000,
         64'h010000008F000000,
         64'h0400000003000000,
         64'h0000000000000000,
         64'h0400000003000000,
         64'h0000000030303030,
         64'h3030634072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h0100000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000000000C00,
         64'h0000000000000002,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0700000001000000,
         64'h0300000001000000,
         64'hC400000010000000,
         64'h0300000000000000,
         64'h30746E696C632C76,
         64'h637369721B000000,
         64'h0D00000003000000,
         64'h0000003030303030,
         64'h303240746E696C63,
         64'h01000000BD000000,
         64'h0000000003000000,
         64'h00007375622D656C,
         64'h706D697300636F73,
         64'h2D657261622D656E,
         64'h616972612C687465,
         64'h1B0000001F000000,
         64'h0300000002000000,
         64'h0F00000004000000,
         64'h0300000002000000,
         64'h0000000004000000,
         64'h0300000000636F73,
         64'h0100000002000000,
         64'h0200000002000000,
         64'h01000000B5000000,
         64'h0400000003000000,
         64'h000063746E692D75,
         64'h70632C7663736972,
         64'h1B0000000F000000,
         64'h03000000A0000000,
         64'h0000000003000000,
         64'h010000008F000000,
         64'h0400000003000000,
         64'h0000000072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h0100000000000000,
         64'h4400000004000000,
         64'h0300000085000000,
         64'h0000000003000000,
         64'h0000393376732C76,
         64'h637369727C000000,
         64'h0B00000003000000,
         64'h00686364616D6966,
         64'h3436767272000000,
         64'h0C00000003000000,
         64'h80F0FA0262000000,
         64'h0400000003000000,
         64'h0000000076637369,
         64'h7200656E61697261,
         64'h2C6874651B000000,
         64'h1100000003000000,
         64'h0000000079616B6F,
         64'h5B00000005000000,
         64'h0300000000757063,
         64'h3800000004000000,
         64'h0300000000000030,
         64'h4075706301000000,
         64'h40787D0148000000,
         64'h0400000003000000,
         64'h000000000F000000,
         64'h0400000003000000,
         64'h0100000000000000,
         64'h0400000003000000,
         64'h0000000073757063,
         64'h0100000002000000,
         64'h0000002000000000,
         64'h0000008000000000,
         64'h4400000010000000,
         64'h0300000000007972,
         64'h6F6D656D38000000,
         64'h0700000003000000,
         64'h0030303030303030,
         64'h384079726F6D656D,
         64'h0100000002000000,
         64'h0000003030323531,
         64'h313A303030303030,
         64'h303440747261752F,
         64'h636F732F2C000000,
         64'h1A00000003000000,
         64'h00006E65736F6863,
         64'h010000000000796D,
         64'h6163636F2C687465,
         64'h260000000B000000,
         64'h0300000000007665,
         64'h642D796D6163636F,
         64'h2C6874651B000000,
         64'h0F00000003000000,
         64'h020000000F000000,
         64'h0400000003000000,
         64'h0200000000000000,
         64'h0400000003000000,
         64'h0000000001000000,
         64'h0000000000000000,
         64'h0000000000000000,
         64'hA805000041010000,
         64'h0000000010000000,
         64'h1100000028000000,
         64'hE005000038000000,
         64'h21070000EDFE0DD0,
         64'h0000001300010020,
         64'hFFDFF06F10500073,
         64'h189000EF9902E283,
         64'h0000129730529073,
         64'h0182829300000297,
         64'hFF8101131BFF8117
    };
    logic [$clog2(RomSize)-1:0] addr_q;
    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end
    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
