/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 713;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h0000000a_0d2e2e2e,
        64'h65646f63_20656874,
        64'h20676e69_74696157,
        64'h00000000_0a0d2164,
        64'h6c726f77_20746f6f,
        64'h62206120_73277449,
        64'h00000000_68746469,
        64'h772d6f69_2d676572,
        64'h00746669_68732d67,
        64'h65720073_74707572,
        64'h7265746e_6900746e,
        64'h65726170_2d747075,
        64'h72726574_6e690064,
        64'h65657073_2d746e65,
        64'h72727563_00766564,
        64'h6e2c7663_73697200,
        64'h79746972_6f697270,
        64'h2d78616d_2c766373,
        64'h69720073_656d616e,
        64'h2d676572_00646564,
        64'h6e657478_652d7374,
        64'h70757272_65746e69,
        64'h00736567_6e617200,
        64'h656c646e_61687000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_00736c6c,
        64'h65632d74_70757272,
        64'h65746e69_23007469,
        64'h6c70732d_626c7400,
        64'h65707974_2d756d6d,
        64'h00617369_2c766373,
        64'h69720073_75746174,
        64'h73006765_72006570,
        64'h79745f65_63697665,
        64'h64007963_6e657571,
        64'h6572662d_6b636f6c,
        64'h63007963_6e657571,
        64'h6572662d_65736162,
        64'h656d6974_00687461,
        64'h702d7475_6f647473,
        64'h006c6564_6f6d0065,
        64'h6c626974_61706d6f,
        64'h6300736c_6c65632d,
        64'h657a6973_2300736c,
        64'h6c65632d_73736572,
        64'h64646123_09000000,
        64'h02000000_02000000,
        64'h02000000_006c6f72,
        64'h746e6f63_d8000000,
        64'h08000000_03000000,
        64'h02000000_0e010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_1f010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h34010000_04000000,
        64'h03000000_02000000,
        64'h2a010000_04000000,
        64'h03000000_01000000,
        64'h1f010000_04000000,
        64'h03000000_02000000,
        64'h0e010000_04000000,
        64'h03000000_80250000,
        64'h00010000_04000000,
        64'h03000000_80969800,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000040,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_d8000000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h01000000_c4000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_f5000000,
        64'h04000000_03000000,
        64'h07000000_e2000000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h01000000_0b000000,
        64'h01000000_c4000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_d8000000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h01000000_03000000,
        64'h01000000_c4000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hbd000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_00000040,
        64'h00000000_00000080,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007972_6f6d656d,
        64'h5b000000_07000000,
        64'h03000000_00303030,
        64'h30303030_38407972,
        64'h6f6d656d_01000000,
        64'h02000000_02000000,
        64'h02000000_01000000,
        64'hb5000000_04000000,
        64'h03000000_00006374,
        64'h6e692d75_70632c76,
        64'h63736972_1b000000,
        64'h0f000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h85000000_00000000,
        64'h03000000_00003933,
        64'h76732c76_63736972,
        64'h7c000000_0b000000,
        64'h03000000_00006364,
        64'h66616d69_34367672,
        64'h72000000_0b000000,
        64'h03000000_00000076,
        64'h63736972_00656e61,
        64'h69726120_2c687465,
        64'h1b000000_12000000,
        64'h03000000_00000000,
        64'h79616b6f_6b000000,
        64'h05000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00757063_5b000000,
        64'h04000000_03000000,
        64'h80969800_4b000000,
        64'h04000000_03000000,
        64'h00000030_40757063,
        64'h01000000_40597307,
        64'h38000000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h73757063_01000000,
        64'h02000000_00303036,
        64'h393a3030_30303030,
        64'h30344074_7261752f,
        64'h636f732f_2c000000,
        64'h18000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hac050000_41010000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'he4050000_38000000,
        64'h25070000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha001ec2f_f0ef8965,
        64'h05130000_15179002,
        64'h16058593_00000597,
        64'hf1402573_edcff0ef,
        64'h89850513_00001517,
        64'hea4ff0ef_e4066805,
        64'h05135805_85931141,
        64'h00989537_6589bba5,
        64'hf00ff0ef_bcc50513,
        64'h00001517_b3dd9265,
        64'h05130000_1517f98f,
        64'hf0ef8526_f1cff0ef,
        64'ha2850513_00001517,
        64'hf28ff0ef_a1c50513,
        64'h00001517_c50d84aa,
        64'hc33ff0ef_9e0d2605,
        64'h8556020a_2583028a,
        64'h3603f4af_f0efbfe5,
        64'h05130000_1517f569,
        64'h93e30804_8493f5ef,
        64'hf0ef2985_97c50513,
        64'h00001517_ff2b9be3,
        64'h835ff0ef_09050009,
        64'h4503f7af_f0efc1e5,
        64'h05130000_1517809f,
        64'hf0ef7088_f8cff0ef,
        64'hc2050513_00001517,
        64'h81bff0ef_6c88f9ef,
        64'hf0efc225_05130000,
        64'h151782df_f0ef0704,
        64'h8b930284_89136888,
        64'hfb8ff0ef_c2c50513,
        64'h00001517_ff2b9be3,
        64'h88dff0ef_09050009,
        64'h45030109_0b93fd6f,
        64'hf0efc2a5_05130000,
        64'h1517fe99_1be38abf,
        64'hf0ef0905_00094503,
        64'hff048913_ff4ff0ef,
        64'hc2850513_00001517,
        64'h8c5ff0ef_0ff9f513,
        64'h809ff0ef_c2450513,
        64'h00001517_b5fda2e5,
        64'h05130000_15178a1f,
        64'hf0ef854e_825ff0ef,
        64'hb3050513_00001517,
        64'h831ff0ef_b2450513,
        64'h00001517_c50d0804,
        64'h89aa8a0a_d3fff0ef,
        64'h850a4605_71010489,
        64'h2583853f_f0efa6e5,
        64'h05130000_15178a1f,
        64'hf0ef4556_865ff0ef,
        64'hc6050513_00001517,
        64'h8b3ff0ef_4546877f,
        64'hf0efc525_05130000,
        64'h1517905f_f0ef6526,
        64'h889ff0ef_c4450513,
        64'h00001517_917ff0ef,
        64'h750289bf_f0efc465,
        64'h05130000_1517929f,
        64'hf0ef6562_8adff0ef,
        64'hc4050513_00001517,
        64'h8fbff0ef_45528bff,
        64'hf0efc425_05130000,
        64'h151790df_f0ef4542,
        64'h8d1ff0ef_c4450513,
        64'h00001517_91fff0ef,
        64'h45328e3f_f0efc465,
        64'h05130000_1517931f,
        64'hf0ef4522_8f5ff0ef,
        64'hc4850513_00001517,
        64'h983ff0ef_4b116502,
        64'h909ff0ef_c4c50513,
        64'h00001517_915ff0ef,
        64'hc3850513_00001517,
        64'hbf6954f9_925ff0ef,
        64'hb4050513_00001517,
        64'h9b3ff0ef_8526937f,
        64'hf0efc425_05130000,
        64'h1517943f_f0efc365,
        64'h05130000_1517c905,
        64'h84aa890a_e4fff0ef,
        64'h850a4585_46057101,
        64'h961ff0ef_c3c50513,
        64'h00001517_80826161,
        64'h6ba26b42_6ae27a02,
        64'h79a27942_74e26406,
        64'h852660a6_fb040113,
        64'h54fd98bf_f0efc3e5,
        64'h05130000_1517c515,
        64'hdf7ff0ef_8aaa0880,
        64'he45ee85a_f052f44e,
        64'hf84afc26_e486ec56,
        64'he0a2715d_b7655479,
        64'h80826169_6baa6b4a,
        64'h6aea7a0a_79aa794a,
        64'h74ea640e_60ae8522,
        64'h547d9d3f_f0efc5e5,
        64'h05130000_1517c59f,
        64'hf0efc5df_f0efc61f,
        64'hf0efc65f_f0efc69f,
        64'hf0efc6df_f0efc71f,
        64'hf0efc75f_f0efa805,
        64'hc7bff0ef_c87ff0ef,
        64'h45314581_46054401,
        64'hf93046e3_19fda17f,
        64'hf0efcc25_05130000,
        64'h1517e799_0359e7b3,
        64'h07241a63_29019041,
        64'h14428c49_cafff0ef,
        64'h90410305_141384a2,
        64'h0085151b_cbfff0ef,
        64'hfd641ae3_04040413,
        64'hff7497e3_892af13f,
        64'hf0ef0485_854a0007,
        64'hc5830094_07b30400,
        64'h0b934481_c67ff0ef,
        64'h850a0400_05938622,
        64'h49018426_20048b13,
        64'hff451ee3_cffff0ef,
        64'h3e800a93_0fe00a13,
        64'he951d15f_f0ef4549,
        64'h85a20ff6_76130016,
        64'h66130015_161bf49f,
        64'hf0ef0ff4_7593f51f,
        64'hf0ef0ff5_f5930084,
        64'h559bf5df_f0ef0ff5,
        64'hf5930104_559bf69f,
        64'hf0ef4501_0ff5f593,
        64'h0184559b_fee79be3,
        64'h078500c6_802300f1,
        64'h06b30800_0713567d,
        64'h47810209_d993842e,
        64'h84aae55e_e95aed56,
        64'hf152f94a_e586fd26,
        64'he1a20206_1993f54e,
        64'h71558082_91411542,
        64'h8d3d8ff9_0057979b,
        64'h17016709_0107d79b,
        64'h0105179b_4105551b,
        64'h0105151b_8d2d00c5,
        64'h95138da9_893d0045,
        64'hd51b8da9_91411542,
        64'h8d5d0522_0085579b,
        64'h808207f5_75138d2d,
        64'h00451593_8d2d8d3d,
        64'h0045d51b_0075d79b,
        64'h8de98082_0141853e,
        64'h640260a2_4781c111,
        64'h57f5f89f_f0efc511,
        64'h57f9efbf_f0efc911,
        64'h57fdeb7f_f0effc6d,
        64'he03ff0ef_347d4429,
        64'hb91ff0ef_e0450513,
        64'h00001517_c89ff0ef,
        64'he022e406_11418082,
        64'h61050015_351364a2,
        64'h644260e2_0004051b,
        64'hfc940ce3_e37ff0ef,
        64'heb3ff0ef_e2c50513,
        64'h00001517_85aa842a,
        64'he53ff0ef_02900513,
        64'h400005b7_07700613,
        64'hfbdff0ef_4485e822,
        64'hec06e426_11018082,
        64'h01410015_3513157d,
        64'h640260a2_0004051b,
        64'hef3ff0ef_e6650513,
        64'h85a20000_1517e89f,
        64'hf0ef842a_e97ff0ef,
        64'he022e406_03700513,
        64'h45810650_06131141,
        64'h80826105_690264a2,
        64'h644260e2_00153513,
        64'hf5650513_0004051b,
        64'h01249863_88bd00f9,
        64'h1b634501_4785ec9f,
        64'hf0efecdf_f0ef842a,
        64'hed3ff0ef_84aaed9f,
        64'hf0efeddf_f0efee1f,
        64'hf0ef892a_eefff0ef,
        64'he04ae426_e822ec06,
        64'h45211aa0_05930870,
        64'h06131101_bfcd4501,
        64'h80826105_690264a2,
        64'h644260e2_4505f89f,
        64'hf0ef4585_ef450513,
        64'h00001517_fe9915e3,
        64'hc00df25f_f0ef892a,
        64'h347df35f_f0ef4501,
        64'h45810950_06134485,
        64'h71040413_e04aec06,
        64'he4266409_e8221101,
        64'hcd1ff06f_6105eee5,
        64'h05130000_151760e2,
        64'h6442da7f_f0ef852e,
        64'h65a2cebf_f0eff365,
        64'h05130000_1517cf7f,
        64'hf0ef8522_cfdff0ef,
        64'he42eec06_f3c50513,
        64'h00001517_842ae822,
        64'h11018082_614564e2,
        64'h740270a2_f47d147d,
        64'h0007d463_4187d79b,
        64'h0185179b_fa7ff0ef,
        64'heb5ff0ef_85320640,
        64'h04136622_ec1ff0ef,
        64'h0ff47513_ec9ff0ef,
        64'h0ff57513_0084551b,
        64'hed5ff0ef_0ff57513,
        64'h0104551b_ee1ff0ef,
        64'h0ff57513_0184551b,
        64'heedff0ef_0404e513,
        64'hfebff0ef_84aa842e,
        64'hec26f022_e432f406,
        64'h7179f07f_f06f0ff0,
        64'h05138082_557db7e9,
        64'h00d70023_078500f6,
        64'h073306c8_2683ff79,
        64'h8b055178_bf4dd6b8,
        64'h07850007_c7038082,
        64'h4501d3b8_4719dbb8,
        64'h577d2000_07b700b6,
        64'hef630007_869b2000,
        64'h08372000_0537fff5,
        64'h8b85537c_20000737,
        64'hd3b82000_07b71060,
        64'h0713fff5_37fd0001,
        64'h03200793_04b76163,
        64'h40a7873b_87aa2000,
        64'h06b7dbb8_57792000,
        64'h07b706b7_ec631000,
        64'h07938082_610564a2,
        64'hd3b84719_dbb86442,
        64'h60e20ff4_7513577d,
        64'h200007b7_e25ff0ef,
        64'h04050513_00001517,
        64'heb3ff0ef_91011502,
        64'h4088e3bf_f0ef05e5,
        64'h05130000_1517e395,
        64'h8b852401_53fc57e0,
        64'hff658b05_06478493,
        64'h53f8d3b8_10600713,
        64'h200007b7_fff537fd,
        64'h00010640_0793d7a8,
        64'hdbb85779_e426e822,
        64'hec062000_07b71101,
        64'he81ff06f_610508e5,
        64'h05130000_151764a2,
        64'h60e26442_d03c4799,
        64'he99ff0ef_0b450513,
        64'h00001517_f27ff0ef,
        64'h91010204_95132481,
        64'heb1ff0ef_0ac50513,
        64'h00001517_5064d03c,
        64'h16600793_ec5ff0ef,
        64'h0e050513_00001517,
        64'hf53ff0ef_91010204,
        64'h95132481_eddff0ef,
        64'h0d850513_00001517,
        64'h5064d03c_10400793,
        64'h20000437_fff537fd,
        64'h000147a9_c3b84729,
        64'h200007b7_f05ff0ef,
        64'he426e822_ec060f85,
        64'h05131101_00001517,
        64'h80824108_8082c10c,
        64'h80826105_60e2ecff,
        64'hf0ef0091_4503ed7f,
        64'hf0ef0081_4503f55f,
        64'hf0efec06_002c1101,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hef9ff0ef_00914503,
        64'hf01ff0ef_34610081,
        64'h4503f81f_f0ef0ff5,
        64'h7513002c_00895533,
        64'h54e10380_0413892a,
        64'hf406e84a_ec26f022,
        64'h71798082_61456942,
        64'h64e27402_70a2fe94,
        64'h10e3f3bf_f0ef0091,
        64'h4503f43f_f0ef3461,
        64'h00814503_fc3ff0ef,
        64'h0ff57513_002c0089,
        64'h553b54e1_4461892a,
        64'hf406e84a_ec26f022,
        64'h71798082_00f58023,
        64'h0007c783_00e580a3,
        64'h97aa8111_00074703,
        64'h973e00f5_771396e7,
        64'h87930000_1797b7f5,
        64'h0405f93f_f0ef8082,
        64'h01416402_60a2e509,
        64'h00044503_842ae406,
        64'he0221141_808200e7,
        64'h88230200_071300e7,
        64'h8423fc70_071300e7,
        64'h8623470d_00a78223,
        64'h0ff57513_00e78023,
        64'h0085551b_0ff57713,
        64'h00e78623_f8000713,
        64'h00078223_400007b7,
        64'h02b5553b_0045959b,
        64'h808200a7_0023dfe5,
        64'h0207f793_01474783,
        64'h40000737_80820205,
        64'h75130147_c5034000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_b8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h25f000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
