package gpio_pkg;

typedef struct packed {
	logic gpio0_d_o;
	logic gpio0_o;
	logic gpio1_d_o;
	logic gpio1_o;
	logic gpio2_d_o;
	logic gpio2_o;
	logic gpio3_d_o;
	logic gpio3_o;
	logic gpio4_d_o;
	logic gpio4_o;
	logic gpio5_d_o;
	logic gpio5_o;
	logic gpio6_d_o;
	logic gpio6_o;
	logic gpio7_d_o;
	logic gpio7_o;
	logic gpio8_d_o;
	logic gpio8_o;
	logic gpio9_d_o;
	logic gpio9_o;
	logic gpio10_d_o;
	logic gpio10_o;
	logic gpio11_d_o;
	logic gpio11_o;
	logic gpio12_d_o;
	logic gpio12_o;
	logic gpio13_d_o;
	logic gpio13_o;
	logic gpio14_d_o;
	logic gpio14_o;
	logic gpio15_d_o;
	logic gpio15_o;
	logic gpio16_d_o;
	logic gpio16_o;
	logic gpio17_d_o;
	logic gpio17_o;
	logic gpio18_d_o;
	logic gpio18_o;
	logic gpio19_d_o;
	logic gpio19_o;
	logic gpio20_d_o;
	logic gpio20_o;
	logic gpio21_d_o;
	logic gpio21_o;
	logic gpio22_d_o;
	logic gpio22_o;
	logic gpio23_d_o;
	logic gpio23_o;
	logic gpio24_d_o;
	logic gpio24_o;
	logic gpio25_d_o;
	logic gpio25_o;
	logic gpio26_d_o;
	logic gpio26_o;
	logic gpio27_d_o;
	logic gpio27_o;
	logic gpio28_d_o;
	logic gpio28_o;
	logic gpio29_d_o;
	logic gpio29_o;
	logic gpio30_d_o;
	logic gpio30_o;
	logic gpio31_d_o;
	logic gpio31_o;
	logic gpio32_d_o;
	logic gpio32_o;
	logic gpio33_d_o;
	logic gpio33_o;
	logic gpio34_d_o;
	logic gpio34_o;
	logic gpio35_d_o;
	logic gpio35_o;
	logic gpio36_d_o;
	logic gpio36_o;
	logic gpio37_d_o;
	logic gpio37_o;
	logic gpio38_d_o;
	logic gpio38_o;
	logic gpio39_d_o;
	logic gpio39_o;
	logic gpio40_d_o;
	logic gpio40_o;
	logic gpio41_d_o;
	logic gpio41_o;
	logic gpio42_d_o;
	logic gpio42_o;
	logic gpio43_d_o;
	logic gpio43_o;
	logic gpio44_d_o;
	logic gpio44_o;
	logic gpio45_d_o;
	logic gpio45_o;
	logic gpio46_d_o;
	logic gpio46_o;
	logic gpio47_d_o;
	logic gpio47_o;
	logic gpio48_d_o;
	logic gpio48_o;
	logic gpio49_d_o;
	logic gpio49_o;
	logic gpio50_d_o;
	logic gpio50_o;
	logic gpio51_d_o;
	logic gpio51_o;
	logic gpio52_d_o;
	logic gpio52_o;
	logic gpio53_d_o;
	logic gpio53_o;
	logic gpio54_d_o;
	logic gpio54_o;
	logic gpio55_d_o;
	logic gpio55_o;
	logic gpio56_d_o;
	logic gpio56_o;
	logic gpio57_d_o;
	logic gpio57_o;
	logic gpio58_d_o;
	logic gpio58_o;
	logic gpio59_d_o;
	logic gpio59_o;
	logic gpio60_d_o;
	logic gpio60_o;
	logic gpio61_d_o;
	logic gpio61_o;
  logic gpio62_d_o;
  logic gpio62_o;
} gpio_to_pad_t;

typedef struct packed {
	logic gpio0_i;
	logic gpio1_i;
	logic gpio2_i;
	logic gpio3_i;
	logic gpio4_i;
	logic gpio5_i;
	logic gpio6_i;
	logic gpio7_i;
	logic gpio8_i;
	logic gpio9_i;
	logic gpio10_i;
	logic gpio11_i;
	logic gpio12_i;
	logic gpio13_i;
	logic gpio14_i;
	logic gpio15_i;
	logic gpio16_i;
	logic gpio17_i;
	logic gpio18_i;
	logic gpio19_i;
	logic gpio20_i;
	logic gpio21_i;
	logic gpio22_i;
	logic gpio23_i;
	logic gpio24_i;
	logic gpio25_i;
	logic gpio26_i;
	logic gpio27_i;
	logic gpio28_i;
	logic gpio29_i;
	logic gpio30_i;
	logic gpio31_i;
	logic gpio32_i;
	logic gpio33_i;
	logic gpio34_i;
	logic gpio35_i;
	logic gpio36_i;
	logic gpio37_i;
	logic gpio38_i;
	logic gpio39_i;
	logic gpio40_i;
	logic gpio41_i;
	logic gpio42_i;
	logic gpio43_i;
	logic gpio44_i;
	logic gpio45_i;
	logic gpio46_i;
	logic gpio47_i;
	logic gpio48_i;
	logic gpio49_i;
	logic gpio50_i;
	logic gpio51_i;
	logic gpio52_i;
	logic gpio53_i;
	logic gpio54_i;
	logic gpio55_i;
	logic gpio56_i;
	logic gpio57_i;
	logic gpio58_i;
	logic gpio59_i;
	logic gpio60_i;
	logic gpio61_i;
  logic gpio62_i;
} pad_to_gpio_t;


endpackage
   
