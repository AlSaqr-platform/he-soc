/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */
// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 301;
    const logic [RomSize-1:0][63:0] mem = {
         64'h4645444342413938,
         64'h3736353433323130,
         64'hFE5FF06F00028067,
         64'h0005628310404537,
         64'h0207A223FEE69CE3,
         64'h0247A68310500073,
         64'h00100713104047B7,
         64'h70858593FFFFF597,
         64'hF140257300008067,
         64'h0201011301813083,
         64'hE65FF0EF00914503,
         64'hE6DFF0EF00814503,
         64'hF09FF0EF00113C23,
         64'h00810593FE010113,
         64'h0000806703010113,
         64'h0101390301813483,
         64'h0201340302813083,
         64'hFC941EE3EA1FF0EF,
         64'h00914503EA9FF0EF,
         64'hFF84041B00814503,
         64'hF49FF0EF0FF57513,
         64'h0081059300895533,
         64'hFF80049303800413,
         64'h0005091302113423,
         64'h0121382300913C23,
         64'h02813023FD010113,
         64'h0000806703010113,
         64'h0101390301813483,
         64'h0201340302813083,
         64'hFC941EE3F01FF0EF,
         64'h00914503F09FF0EF,
         64'hFF84041B00814503,
         64'hFA9FF0EF0FF57513,
         64'h008105930089553B,
         64'hFF80049301800413,
         64'h0005091302113423,
         64'h0121382300913C23,
         64'h02813023FD010113,
         64'h0000806700F58023,
         64'h0007C78300E580A3,
         64'h00A787B300455513,
         64'h0007470300E78733,
         64'h00F5771314C78793,
         64'h00000797FE1FF06F,
         64'h00140413F79FF0EF,
         64'h0000806701010113,
         64'h0001340300813083,
         64'h00051A6300044503,
         64'h0005041300113423,
         64'h00813023FF010113,
         64'h0000806700E78823,
         64'h0200071300E78423,
         64'hFC70071300E78623,
         64'h0030071300A78223,
         64'h0FF5751300E78023,
         64'h0085551B0FF57713,
         64'h00E78623F8000713,
         64'h00078223400007B7,
         64'h02B5553B0045959B,
         64'h0000806700A70023,
         64'hFE078CE30207F793,
         64'h0147478340000737,
         64'h0000806702057513,
         64'h0147C503400007B7,
         64'h0000806700054503,
         64'h0000806700B50023,
         64'h0000806700000000,
         64'h68746469772D6F69,
         64'h2D67657200746669,
         64'h68732D6765720073,
         64'h747075727265746E,
         64'h6900746E65726170,
         64'h2D74707572726574,
         64'h6E69006465657073,
         64'h2D746E6572727563,
         64'h007665646E2C7663,
         64'h7369720079746972,
         64'h6F6972702D78616D,
         64'h2C76637369720073,
         64'h656D616E2D676572,
         64'h006465646E657478,
         64'h652D737470757272,
         64'h65746E6900736567,
         64'h6E617200656C646E,
         64'h6168700072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h00736C6C65632D74,
         64'h7075727265746E69,
         64'h230074696C70732D,
         64'h626C740065707974,
         64'h2D756D6D00617369,
         64'h2C76637369720079,
         64'h636E657571657266,
         64'h2D6B636F6C630073,
         64'h7574617473007963,
         64'h6E6575716572662D,
         64'h65736162656D6974,
         64'h0067657200657079,
         64'h745F656369766564,
         64'h00687461702D7475,
         64'h6F647473006C6564,
         64'h6F6D00656C626974,
         64'h61706D6F6300736C,
         64'h6C65632D657A6973,
         64'h2300736C6C65632D,
         64'h7373657264646123,
         64'h0900000002000000,
         64'h0200000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000002000000,
         64'h0E01000004000000,
         64'h0300000000100000,
         64'h0000000000000018,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0700000006000000,
         64'h0500000004000000,
         64'h1F01000010000000,
         64'h0300000000007265,
         64'h6D69745F6270612C,
         64'h706C75701B000000,
         64'h0F00000003000000,
         64'h0000303030303030,
         64'h38314072656D6974,
         64'h0100000002000000,
         64'h0400000034010000,
         64'h0400000003000000,
         64'h020000002A010000,
         64'h0400000003000000,
         64'h020000001F010000,
         64'h0400000003000000,
         64'h020000000E010000,
         64'h0400000003000000,
         64'h00C2010000010000,
         64'h0400000003000000,
         64'h80F0FA0262000000,
         64'h0400000003000000,
         64'h0010000000000000,
         64'h0000004000000000,
         64'h4400000010000000,
         64'h0300000000303535,
         64'h3631736E1B000000,
         64'h0800000003000000,
         64'h0000003030303030,
         64'h3030344074726175,
         64'h0100000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000000100000,
         64'h0000000000000000,
         64'h0000000044000000,
         64'h1000000003000000,
         64'hFFFF000001000000,
         64'hC400000008000000,
         64'h0300000000333130,
         64'h2D67756265642C76,
         64'h637369721B000000,
         64'h1000000003000000,
         64'h0000304072656C6C,
         64'h6F72746E6F632D67,
         64'h7562656401000000,
         64'h0200000002000000,
         64'hB500000004000000,
         64'h03000000FF000000,
         64'hF500000004000000,
         64'h0300000007000000,
         64'hE200000004000000,
         64'h0300000000000004,
         64'h000000000000000C,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0900000001000000,
         64'h0B00000001000000,
         64'hC400000010000000,
         64'h03000000A0000000,
         64'h0000000003000000,
         64'h003063696C702C76,
         64'h637369721B000000,
         64'h0C00000003000000,
         64'h010000008F000000,
         64'h0400000003000000,
         64'h0000000000000000,
         64'h0400000003000000,
         64'h0000000030303030,
         64'h3030634072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h0100000002000000,
         64'h006C6F72746E6F63,
         64'hD800000008000000,
         64'h0300000000000C00,
         64'h0000000000000002,
         64'h0000000044000000,
         64'h1000000003000000,
         64'h0700000001000000,
         64'h0300000001000000,
         64'hC400000010000000,
         64'h0300000000000000,
         64'h30746E696C632C76,
         64'h637369721B000000,
         64'h0D00000003000000,
         64'h0000003030303030,
         64'h303240746E696C63,
         64'h01000000BD000000,
         64'h0000000003000000,
         64'h00007375622D656C,
         64'h706D697300636F73,
         64'h2D657261622D656E,
         64'h616972612C687465,
         64'h1B0000001F000000,
         64'h0300000002000000,
         64'h0F00000004000000,
         64'h0300000002000000,
         64'h0000000004000000,
         64'h0300000000636F73,
         64'h0100000002000000,
         64'h0200000002000000,
         64'h01000000B5000000,
         64'h0400000003000000,
         64'h000063746E692D75,
         64'h70632C7663736972,
         64'h1B0000000F000000,
         64'h03000000A0000000,
         64'h0000000003000000,
         64'h010000008F000000,
         64'h0400000003000000,
         64'h0000000072656C6C,
         64'h6F72746E6F632D74,
         64'h7075727265746E69,
         64'h0100000000000000,
         64'h4400000004000000,
         64'h0300000085000000,
         64'h0000000003000000,
         64'h0000393376732C76,
         64'h637369727C000000,
         64'h0B00000003000000,
         64'h00686364616D6966,
         64'h3436767272000000,
         64'h0C00000003000000,
         64'h80F0FA0262000000,
         64'h0400000003000000,
         64'h0000000076637369,
         64'h7200656E61697261,
         64'h2C6874651B000000,
         64'h1100000003000000,
         64'h0000000079616B6F,
         64'h5B00000005000000,
         64'h0300000000757063,
         64'h3800000004000000,
         64'h0300000000000030,
         64'h4075706301000000,
         64'h40787D0148000000,
         64'h0400000003000000,
         64'h000000000F000000,
         64'h0400000003000000,
         64'h0100000000000000,
         64'h0400000003000000,
         64'h0000000073757063,
         64'h0100000002000000,
         64'h0000002000000000,
         64'h0000008000000000,
         64'h4400000010000000,
         64'h0300000000007972,
         64'h6F6D656D38000000,
         64'h0700000003000000,
         64'h0030303030303030,
         64'h384079726F6D656D,
         64'h0100000002000000,
         64'h0000003030323531,
         64'h313A303030303030,
         64'h303440747261752F,
         64'h636F732F2C000000,
         64'h1A00000003000000,
         64'h00006E65736F6863,
         64'h010000000000796D,
         64'h6163636F2C687465,
         64'h260000000B000000,
         64'h0300000000007665,
         64'h642D796D6163636F,
         64'h2C6874651B000000,
         64'h0F00000003000000,
         64'h020000000F000000,
         64'h0400000003000000,
         64'h0200000000000000,
         64'h0400000003000000,
         64'h0000000001000000,
         64'h0000000000000000,
         64'h0000000000000000,
         64'hA805000041010000,
         64'h0000000010000000,
         64'h1100000028000000,
         64'hE005000038000000,
         64'h21070000EDFE0DD0,
         64'h0000001300010020,
         64'hFFDFF06F10500073,
         64'h109000EF9102E283,
         64'h0000129730529073,
         64'h0182829300000297,
         64'h01A111130210011B
    };
    logic [$clog2(RomSize)-1:0] addr_q;
    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end
    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
